
class zuspec_component;
endclass
