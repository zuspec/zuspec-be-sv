
package zuspec;

endpackage

